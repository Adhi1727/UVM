VSIMSA: Configuration file changed: `/home/runner/library.cfg'
ALIB: Library "work" attached.
work = ./work/work.lib
MESSAGE_SP VCP2124 "Package uvm_pkg found in library uvm_1_2."
MESSAGE "Unit top modules: top."
SUCCESS "Compile success 0 Errors 0 Warnings  Analysis time: 5[s]."
done
# Aldec, Inc. Riviera-PRO version 2025.04.139.9738 built for Linux64 on May 30, 2025.
# HDL, SystemC, and Assertions simulator, debugger, and design environment.
# (c) 1999-2025 Aldec, Inc. All rights reserved.
# ELBREAD: Elaboration process.
# ELBREAD: Warning: ELBREAD_0049 The "uvm_pkg" design unit does not have a time unit/precision defined but other design units do.
# ELBREAD: Elaboration time 0.6 [s].
# KERNEL: Main thread initiated.
# KERNEL: Kernel process initialization phase.
# ELAB2: Elaboration final pass...
# KERNEL: PLI/VHPI kernel's engine initialization done.
# PLI: Loading library '/usr/share/Riviera-PRO/bin/libsystf.so'
# ELAB2: Create instances ...
# KERNEL: Info: Loading library:  /usr/share/Riviera-PRO/bin/uvm_1_2_dpi
# KERNEL: Time resolution set to 1ns.
# ELAB2: Create instances complete.
# SLP: Started
# SLP: Elaboration phase ...
# SLP: Elaboration phase ... done : 0.0 [s]
# SLP: Generation phase ...
# SLP: Generation phase ... done : 0.0 [s]
# SLP: Finished : 0.1 [s]
# SLP: 0 primitives and 2 (28.57%) other processes in SLP
# SLP: 20 (0.07%) signals in SLP and 10 (0.03%) interface signals
# ELAB2: Elaboration final pass complete - time: 2.0 [s].
# KERNEL: SLP loading done - time: 0.0 [s].
# KERNEL: Warning: You are using the Riviera-PRO EDU Edition. The performance of simulation is reduced.
# KERNEL: Warning: Contact Aldec for available upgrade options - sales@aldec.com.
# KERNEL: SLP simulation initialization done - time: 0.0 [s].
# KERNEL: Kernel process initialization done.
# Allocation: Simulator allocated 28384 kB (elbread=2094 elab2=21540 kernel=4749 sdf=0)
# KERNEL: UVM_INFO ./uvm-1.2/src/base/uvm_root.svh(392) @ 0: reporter [UVM/RELNOTES] 
# KERNEL: ----------------------------------------------------------------
# KERNEL: UVM-1.2
# KERNEL: (C) 2007-2014 Mentor Graphics Corporation
# KERNEL: (C) 2007-2014 Cadence Design Systems, Inc.
# KERNEL: (C) 2006-2014 Synopsys, Inc.
# KERNEL: (C) 2011-2013 Cypress Semiconductor Corp.
# KERNEL: (C) 2013-2014 NVIDIA Corporation
# KERNEL: ----------------------------------------------------------------
# KERNEL: 
# KERNEL:   ***********       IMPORTANT RELEASE NOTES         ************
# KERNEL: 
# KERNEL:   You are using a version of the UVM library that has been compiled
# KERNEL:   with `UVM_NO_DEPRECATED undefined.
# KERNEL:   See http://www.eda.org/svdb/view.php?id=3313 for more details.
# KERNEL: 
# KERNEL:   You are using a version of the UVM library that has been compiled
# KERNEL:   with `UVM_OBJECT_DO_NOT_NEED_CONSTRUCTOR undefined.
# KERNEL:   See http://www.eda.org/svdb/view.php?id=3770 for more details.
# KERNEL: 
# KERNEL:       (Specify +UVM_NO_RELNOTES to turn off this notice)
# KERNEL: 
# KERNEL: ASDB file was created in location /home/runner/dataset.asdb
# KERNEL: UVM_INFO @ 0: reporter [RNTST] Running test test...
# KERNEL: UVM_INFO /home/runner/env.sv(10) @ 0: uvm_test_top.en [ENV] environment created
# KERNEL: UVM_INFO /home/runner/fa_sequencer.sv(8) @ 0: uvm_test_top.en.agn.seqr [SEQ_R] Sequencer created
# KERNEL: UVM_INFO /home/runner/fa_sequence.sv(12) @ 0: uvm_test_top.en.agn.seqr@@se [SEQ] sequence started
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 10: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 20: uvm_test_top.en.score [SCAD] PASS! input: a = 0 | b = 1 | cin = 1 output: sum = 0 | cout = 1
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 30: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 40: uvm_test_top.en.score [SCAD] PASS! input: a = 0 | b = 1 | cin = 1 output: sum = 0 | cout = 1
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 50: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 60: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 70: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 80: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# KERNEL: UVM_INFO /home/runner/scoreboard.sv(25) @ 90: uvm_test_top.en.score [SCAD] PASS! input: a = 1 | b = 0 | cin = 0 output: sum = 1 | cout = 0
# RUNTIME: Info: RUNTIME_0068 testbench.sv (36): $finish called.
# KERNEL: Time: 100 ns,  Iteration: 0,  Instance: /top,  Process: @INITIAL#32_1@.
# KERNEL: stopped at time: 100 ns
# VSIM: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
