interface dff_interface;
  logic clk;
  logic rst;
  logic d;
  logic q;
endinterface
