interface fa_interface;
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic cout;
endinterface
