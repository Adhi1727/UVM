You are using a version of the UVM library that has been compiled
  with `UVM_NO_DEPRECATED undefined.
  See http://www.eda.org/svdb/view.php?id=3313 for more details.

  You are using a version of the UVM library that has been compiled
  with `UVM_OBJECT_DO_NOT_NEED_CONSTRUCTOR undefined.
  See http://www.eda.org/svdb/view.php?id=3770 for more details.

      (Specify +UVM_NO_RELNOTES to turn off this notice)

UVM_INFO @ 0: reporter [RNTST] Running test test...
UVM_INFO sequencer.sv(6) @ 0: uvm_test_top.en.agnt.seqr [SEQR] Sequencer Created
UVM_INFO sequence.sv(11) @ 0: uvm_test_top.en.agnt.seqr@@seq [SEQ] Sequence Started
UVM_INFO scoreboard.sv(25) @ 6: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 16: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 26: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 36: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 46: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 56: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 66: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 76: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 86: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 96: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 106: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 116: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 126: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 136: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 146: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 156: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=1|Actual output: q=1|| Expected output: q=1
UVM_INFO scoreboard.sv(25) @ 166: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=0|d=1|Actual output: q=1|| Expected output: q=1
UVM_INFO scoreboard.sv(25) @ 176: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 186: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 196: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 206: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 216: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 226: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 236: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 246: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 256: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 266: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 276: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 286: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
UVM_INFO scoreboard.sv(25) @ 296: uvm_test_top.en.score [SB] PASS----> INPUT:clk=0 |rst=1|d=0|Actual output: q=0|| Expected output: q=0
$finish called from file "testbench.sv", line 36.
$finish at simulation time                  300
           V C S   S i m u l a t i o n   R e p o r t 
Time: 300 ns
CPU Time:      0.640 seconds;  
